/* verilator lint_off UNPACKED */
/* verilator lint_off WIDTH */
/* verilator lint_off UNUSED */
/* verilator lint_off UNDRIVEN */

module memory 
#( 
	parameter data_width 	= 8,
	parameter weight_width 	= 8
) (	
	input logic clk,
	input logic rstn,
	
	input logic	     mode,
	input logic [31 : 0] data_idx,
	input logic [31 : 0] weight_idx,
	input logic [31 : 0] result_idx,
	input logic	     write_enable,

	input logic  [  data_width-1 : 0] result,
	output logic [  data_width-1 : 0] data,
	output logic [weight_width-1 : 0] weight
);


    logic [  data_width-1 : 0] data_a0, data_a1;

	logic [  data_width-1 : 0] memory_A0 [8191 : 0];
	logic [  data_width-1 : 0] memory_A1 [8191 : 0];
	logic [weight_width-1 : 0] memory_B  [3438-1 : 0] = '{8'b00000000,8'b11110100,8'b00101010,8'b00100101,8'b11101101,8'b00001101,8'b00000010,8'b00000011,8'b11011111,8'b00011101,8'b11100011,8'b00011000,8'b00001001,8'b00000000,8'b00000110,8'b11111001,8'b00001111,8'b11101001,8'b00000101,8'b11111110,8'b11110111,8'b00010100,8'b11110111,8'b11110001,8'b00011010,8'b11010100,8'b00001011,8'b11011100,8'b00001001,8'b00001000,8'b11111010,8'b11111010,8'b11101100,8'b11111100,8'b11011011,8'b11110100,8'b11110111,8'b00000111,8'b11111111,8'b00000101,8'b11101110,8'b00010010,8'b11101001,8'b00011011,8'b00011011,8'b11110000,8'b11110000,8'b00100100,8'b00000101,8'b11110100,8'b00010111,8'b11111001,8'b11111001,8'b00010110,8'b00010010,8'b11111010,8'b11101000,8'b00001101,8'b11001110,8'b00000001,8'b00010010,8'b11110011,8'b11101111,8'b00010010,8'b00001010,8'b11111001,8'b00000010,8'b11111010,8'b11011011,8'b00001110,8'b11110101,8'b11101001,8'b11100101,8'b00001011,8'b10110010,8'b00010100,8'b00000111,8'b11101111,8'b11100110,8'b00001110,8'b00001001,8'b11110011,8'b11100111,8'b00010100,8'b11011000,8'b00010011,8'b11001011,8'b11011010,8'b11011000,8'b00010001,8'b11010011,8'b00001101,8'b00010001,8'b11111111,8'b11101101,8'b00011001,8'b00100001,8'b11101000,8'b00001001,8'b11110111,8'b11110001,8'b00001111,8'b11101111,8'b00000011,8'b11111011,8'b00001011,8'b11011001,8'b00000011,8'b11101010,8'b11111111,8'b00001010,8'b00001101,8'b00000000,8'b11110111,8'b00101101,8'b11111001,8'b11011000,8'b00000011,8'b11011000,8'b11111000,8'b11110010,8'b11110100,8'b11101110,8'b11111101,8'b00001011,8'b00001010,8'b00001010,8'b00000110,8'b00100101,8'b11110011,8'b00001011,8'b11100010,8'b11101010,8'b00010111,8'b11111010,8'b11100101,8'b11011101,8'b00001100,8'b11100110,8'b00000101,8'b11100100,8'b00001001,8'b00110100,8'b11111110,8'b00100000,8'b11110111,8'b00000000,8'b00000111,8'b11111001,8'b00010000,8'b11011010,8'b11101100,8'b11111011,8'b11111111,8'b11011011,8'b00001011,8'b00001000,8'b11111100,8'b00010001,8'b11111011,8'b00010000,8'b11110000,8'b11001110,8'b00001000,8'b11101100,8'b00001011,8'b11110110,8'b11111001,8'b11110010,8'b00001111,8'b00001000,8'b00000100,8'b00000011,8'b11111010,8'b00100001,8'b00001001,8'b00001011,8'b11110001,8'b11110010,8'b11101011,8'b11101100,8'b00010110,8'b11110101,8'b11110000,8'b00001001,8'b11110111,8'b00000110,8'b11001100,8'b11011111,8'b00000110,8'b00000000,8'b11110110,8'b11110111,8'b11110110,8'b00010100,8'b11110111,8'b11110001,8'b11111101,8'b11100010,8'b11111011,8'b00101011,8'b11111110,8'b11011100,8'b11100000,8'b00011111,8'b11110000,8'b11111000,8'b11001000,8'b11010110,8'b00001110,8'b00010001,8'b00001110,8'b11011101,8'b11110010,8'b00100101,8'b11101010,8'b11010001,8'b11110101,8'b11011100,8'b00010111,8'b11111000,8'b11110011,8'b11110010,8'b11110011,8'b00101011,8'b11010010,8'b11110000,8'b10110111,8'b11100110,8'b00001101,8'b11101101,8'b11011011,8'b11101110,8'b00000111,8'b00101100,8'b10111101,8'b11011111,8'b10110110,8'b11100011,8'b00010000,8'b11110000,8'b11010001,8'b11110111,8'b00000001,8'b00010100,8'b10111100,8'b11110111,8'b10001111,8'b11001001,8'b00000111,8'b11101011,8'b11000100,8'b11101000,8'b00001001,8'b00011110,8'b11110100,8'b11111000,8'b11011110,8'b11011101,8'b11111110,8'b11100110,8'b11010010,8'b11110100,8'b00000110,8'b00100111,8'b10110011,8'b00000111,8'b11011011,8'b11010100,8'b11110101,8'b11110110,8'b11001010,8'b11111000,8'b00001011,8'b00100110,8'b11000001,8'b11111000,8'b11001000,8'b11110000,8'b11111101,8'b00000011,8'b11111001,8'b00001101,8'b00000101,8'b00001000,8'b11100100,8'b11110011,8'b11101111,8'b11100100,8'b11100101,8'b00001010,8'b00000001,8'b00000100,8'b00000101,8'b00010110,8'b00001011,8'b11111001,8'b11011101,8'b11110100,8'b00000100,8'b11111111,8'b11111010,8'b00000011,8'b11111010,8'b00001111,8'b00000100,8'b11111000,8'b11001111,8'b00000000,8'b00001000,8'b11111111,8'b11011010,8'b00010001,8'b00000000,8'b00010000,8'b11010101,8'b00000010,8'b11101011,8'b11111110,8'b00010100,8'b11111110,8'b11100111,8'b00001111,8'b00000001,8'b00010010,8'b11010001,8'b00001010,8'b11001110,8'b11110111,8'b00001010,8'b11111110,8'b00000001,8'b00001000,8'b11111001,8'b00001011,8'b11110000,8'b11111101,8'b11010100,8'b11110101,8'b00001011,8'b11111100,8'b00000101,8'b00000101,8'b11111011,8'b00001000,8'b11111001,8'b11111111,8'b11011010,8'b11111010,8'b00000111,8'b00000011,8'b00000000,8'b00001101,8'b00000010,8'b00000011,8'b11110000,8'b11111100,8'b11100001,8'b11110001,8'b00001011,8'b11111111,8'b11110000,8'b00010010,8'b00000001,8'b00000000,8'b11011110,8'b11111111,8'b11010011,8'b11111011,8'b11111101,8'b00000001,8'b00000011,8'b11111010,8'b11111100,8'b00000110,8'b00000001,8'b11111111,8'b00000001,8'b11111000,8'b11100100,8'b11111101,8'b11101111,8'b00000101,8'b00000010,8'b00001001,8'b11111010,8'b00000000,8'b11111101,8'b00001000,8'b11100111,8'b00000000,8'b11101111,8'b00010010,8'b00001100,8'b00010011,8'b11111100,8'b00000101,8'b00001000,8'b00000010,8'b11111000,8'b11111001,8'b11100011,8'b00001101,8'b00000100,8'b00001000,8'b11110011,8'b00000011,8'b00000111,8'b00000001,8'b00000010,8'b11111001,8'b11111111,8'b00001011,8'b11111011,8'b00000111,8'b11100110,8'b11111100,8'b00000000,8'b11110110,8'b00000100,8'b00000010,8'b00001011,8'b00001000,8'b11101000,8'b00000001,8'b11111111,8'b11111110,8'b11111110,8'b11110110,8'b00000101,8'b00000100,8'b00000111,8'b00001001,8'b11001110,8'b11101110,8'b00000010,8'b00000100,8'b00000001,8'b11111110,8'b00000000,8'b00001001,8'b00000111,8'b00000110,8'b11100010,8'b11100000,8'b00000110,8'b00001001,8'b11111110,8'b11111111,8'b00000100,8'b00000100,8'b11111100,8'b00000011,8'b11100101,8'b11101011,8'b11111011,8'b00000001,8'b11110101,8'b00001100,8'b00000101,8'b11101110,8'b11110011,8'b11110110,8'b11111001,8'b00000110,8'b00000000,8'b11111010,8'b00001000,8'b00001000,8'b11011111,8'b11101110,8'b11110000,8'b00000011,8'b00000011,8'b00010101,8'b00000011,8'b00000011,8'b00001011,8'b00000100,8'b11010111,8'b11100110,8'b11101001,8'b00000111,8'b00000011,8'b00000101,8'b00000010,8'b00000001,8'b00000110,8'b00000101,8'b11111000,8'b11101101,8'b11101001,8'b00000110,8'b00000000,8'b00000100,8'b00000000,8'b11111010,8'b11111110,8'b00000011,8'b00000001,8'b11111011,8'b11111101,8'b00000100,8'b11111100,8'b00000100,8'b11110110,8'b11111011,8'b11111011,8'b11111100,8'b00000111,8'b00000110,8'b00001000,8'b00000111,8'b11100101,8'b11111001,8'b00001010,8'b00000111,8'b00001000,8'b00000110,8'b00000100,8'b00001011,8'b00000100,8'b00001010,8'b10110110,8'b11011001,8'b00001001,8'b00000111,8'b00000100,8'b00001010,8'b11111110,8'b00001010,8'b00000010,8'b00000111,8'b10100110,8'b11100110,8'b00000111,8'b00000101,8'b00000011,8'b00001011,8'b11111101,8'b00000111,8'b11111010,8'b00000110,8'b10110011,8'b11111011,8'b00000110,8'b00001110,8'b00000101,8'b00010001,8'b11111111,8'b11110000,8'b11100101,8'b00000010,8'b11101111,8'b00010011,8'b00000110,8'b11110100,8'b00000111,8'b00001001,8'b11110010,8'b11010111,8'b11100111,8'b00001000,8'b11110101,8'b00001100,8'b00000100,8'b11110100,8'b00001001,8'b00001000,8'b11101100,8'b11011111,8'b11110110,8'b00001001,8'b11111110,8'b00001010,8'b00001100,8'b11111100,8'b00001100,8'b00001010,8'b11111010,8'b11110100,8'b11100100,8'b00000110,8'b00000001,8'b00001001,8'b00000010,8'b00000000,8'b11111110,8'b11111100,8'b00000010,8'b00000001,8'b11110011,8'b11110100,8'b11110100,8'b11111111,8'b00000001,8'b00000001,8'b11110010,8'b11111100,8'b00000011,8'b00000101,8'b11110111,8'b00000100,8'b11101111,8'b11110011,8'b00000011,8'b11111111,8'b00000001,8'b00000101,8'b11111110,8'b00000100,8'b11110110,8'b00000010,8'b11110001,8'b11110011,8'b00000101,8'b11111001,8'b11111111,8'b00001001,8'b11110001,8'b00000100,8'b11110010,8'b00000011,8'b11101100,8'b11111111,8'b00000110,8'b11110101,8'b00000000,8'b00001101,8'b11110100,8'b00000011,8'b11101101,8'b00000010,8'b11100100,8'b00000110,8'b00001011,8'b11111001,8'b00000101,8'b00001111,8'b10110110,8'b00001110,8'b11100100,8'b00001000,8'b11101110,8'b00000111,8'b00000100,8'b11101101,8'b11111010,8'b00001111,8'b11011000,8'b00000101,8'b11100011,8'b00000111,8'b11100110,8'b00000111,8'b00000101,8'b11111100,8'b00001011,8'b00001110,8'b11111011,8'b11111110,8'b11010011,8'b00001010,8'b11101011,8'b00001001,8'b00001001,8'b00000011,8'b00000001,8'b00010100,8'b00000111,8'b00001000,8'b11011000,8'b11111111,8'b11110100,8'b00001111,8'b00000010,8'b00010001,8'b11011110,8'b11111010,8'b00000100,8'b00000000,8'b11100101,8'b11111000,8'b11111011,8'b00000101,8'b00000000,8'b00000010,8'b11111101,8'b11111111,8'b00000010,8'b11111111,8'b11111001,8'b11111110,8'b11111101,8'b00000010,8'b00000000,8'b11110110,8'b00000001,8'b00000011,8'b00000000,8'b11111110,8'b00000100,8'b00000000,8'b11111111,8'b00000010,8'b00000100,8'b11110101,8'b00000101,8'b00000101,8'b11001100,8'b11111001,8'b11111111,8'b11111110,8'b11111101,8'b00000001,8'b00001000,8'b11110101,8'b00000101,8'b00001001,8'b11100110,8'b11110100,8'b11111001,8'b11111100,8'b11111010,8'b00000011,8'b00001111,8'b11110011,8'b11111011,8'b00001010,8'b11110001,8'b00001111,8'b11110101,8'b11110111,8'b00000000,8'b11111110,8'b11101011,8'b11111100,8'b11110001,8'b00001011,8'b11111001,8'b00001011,8'b11101001,8'b11101101,8'b11101110,8'b00001001,8'b11111011,8'b00001100,8'b11110010,8'b00010100,8'b00000001,8'b00001111,8'b11100001,8'b11110111,8'b11101101,8'b00010000,8'b11111010,8'b00010000,8'b11011110,8'b00000111,8'b00000101,8'b00000101,8'b11001011,8'b00000000,8'b11110000,8'b00000111,8'b00000011,8'b00001000,8'b11111011,8'b11110110,8'b11111111,8'b11111011,8'b11110101,8'b11111111,8'b11111110,8'b11111010,8'b00000010,8'b11111111,8'b00000011,8'b11111111,8'b11111100,8'b11110111,8'b00000101,8'b00000011,8'b00000011,8'b00000001,8'b00000011,8'b00000010,8'b00000101,8'b00000011,8'b11100111,8'b11111000,8'b00000110,8'b00000010,8'b00000110,8'b00000010,8'b00000100,8'b00000010,8'b00000101,8'b00000001,8'b11100010,8'b11110101,8'b00000100,8'b11111100,8'b00000000,8'b00000001,8'b00000001,8'b11111101,8'b00000010,8'b00001001,8'b11101101,8'b11110100,8'b11111110,8'b11111011,8'b00000101,8'b11111100,8'b00000100,8'b00000100,8'b11111101,8'b00000111,8'b00001110,8'b00000101,8'b00000100,8'b11011010,8'b11111011,8'b11100100,8'b11110001,8'b00000111,8'b11011101,8'b00001000,8'b00001100,8'b00001001,8'b00000000,8'b11101010,8'b00000000,8'b11101010,8'b11110111,8'b00001010,8'b11110100,8'b00001000,8'b00001100,8'b11111110,8'b11100011,8'b00000001,8'b11101100,8'b11111010,8'b00000111,8'b00001100,8'b00000111,8'b11110110,8'b00001011,8'b11101101,8'b11011100,8'b00000100,8'b11110001,8'b11100111,8'b00000111,8'b00000001,8'b00000110,8'b11110110,8'b11111111,8'b11101110,8'b11111010,8'b00000010,8'b00000000,8'b11100011,8'b00000001,8'b00000000,8'b00000011,8'b00000001,8'b11111001,8'b11110000,8'b00000100,8'b00000010,8'b00000100,8'b11111000,8'b00000001,8'b00000101,8'b00000011,8'b00000111,8'b11110101,8'b11110011,8'b00000110,8'b00000000,8'b00000110,8'b11111111,8'b00000001,8'b00000011,8'b00000001,8'b11111110,8'b11111110,8'b11110100,8'b00000110,8'b11110100,8'b00000101,8'b11111100,8'b11111100,8'b00000100,8'b11111110,8'b00001000,8'b00000111,8'b11111010,8'b00000101,8'b11111101,8'b00001101,8'b11101101,8'b11111100,8'b00000100,8'b00000011,8'b11111010,8'b00001110,8'b11101110,8'b00010001,8'b00000010,8'b00000010,8'b10101110,8'b00010101,8'b11110100,8'b00000100,8'b11100110,8'b00001111,8'b11011110,8'b00010011,8'b00000010,8'b00000111,8'b11010011,8'b00011001,8'b11111000,8'b00001001,8'b11011110,8'b00001001,8'b11001000,8'b11110010,8'b00001100,8'b11110010,8'b11000111,8'b00010111,8'b11101011,8'b00010101,8'b10100111,8'b00001011,8'b10100001,8'b11100011,8'b00010110,8'b11101100,8'b11100011,8'b00011011,8'b11101110,8'b00011101,8'b10101010,8'b00001000,8'b10110000,8'b00001000,8'b00010001,8'b00000000,8'b11010000,8'b00010100,8'b11101011,8'b00010101,8'b11001001,8'b00000110,8'b11000011,8'b00001000,8'b00001010,8'b00001000,8'b11001110,8'b00001111,8'b00000010,8'b00001100,8'b11100111,8'b00001010,8'b11100101,8'b00001011,8'b00000011,8'b00001000,8'b11110010,8'b00001011,8'b00000110,8'b00000110,8'b11101000,8'b00000111,8'b11111001,8'b00000110,8'b00000011,8'b00000000,8'b11101000,8'b00000100,8'b11111110,8'b00000011,8'b11011111,8'b00001001,8'b11101110,8'b11101010,8'b00000000,8'b00000111,8'b11100010,8'b11101101,8'b11111010,8'b00010011,8'b11110100,8'b00001000,8'b11100000,8'b00011001,8'b00010000,8'b11100011,8'b00001100,8'b11111101,8'b11011010,8'b11011101,8'b11110000,8'b00010100,8'b00000011,8'b11111100,8'b00001110,8'b11011111,8'b11111110,8'b11110111,8'b11101101,8'b11000010,8'b11111111,8'b00000001,8'b00010101,8'b00001101,8'b00001000,8'b11101111,8'b11110011,8'b11111001,8'b11100110,8'b11001100,8'b11111001,8'b11110110,8'b00001111,8'b00001000,8'b11110000,8'b11101101,8'b11100010,8'b11111000,8'b11110100,8'b11110110,8'b11110010,8'b11110011,8'b00001011,8'b00001001,8'b11010011,8'b11110011,8'b11101001,8'b11101010,8'b11111100,8'b11111110,8'b11111110,8'b11101011,8'b00001110,8'b00000111,8'b11010110,8'b00000001,8'b11111011,8'b11101010,8'b00000101,8'b00000010,8'b11111000,8'b11111110,8'b00000110,8'b00000010,8'b11100100,8'b00000001,8'b00000000,8'b11011010,8'b00000110,8'b00000000,8'b00000000,8'b00000111,8'b00001001,8'b11111011,8'b00000000,8'b00000101,8'b00010100,8'b11000100,8'b00001000,8'b11111010,8'b11110111,8'b00001110,8'b11101110,8'b11100000,8'b00101100,8'b00010000,8'b00011011,8'b11000000,8'b00000110,8'b10110000,8'b11111100,8'b00000110,8'b00000010,8'b00010000,8'b11110110,8'b11001011,8'b00001100,8'b00010000,8'b11010101,8'b10110011,8'b11101011,8'b11111010,8'b00000011,8'b00001011,8'b00000101,8'b11101111,8'b11110101,8'b00010010,8'b11101100,8'b10110101,8'b11110000,8'b11110110,8'b00001011,8'b00001011,8'b11110110,8'b11111100,8'b11100101,8'b00010011,8'b11111101,8'b11101001,8'b11110111,8'b11111001,8'b00000111,8'b00001010,8'b11101011,8'b11111110,8'b11100000,8'b00001101,8'b00000001,8'b11111101,8'b11111100,8'b11110001,8'b00000111,8'b00000110,8'b11001111,8'b00000100,8'b11101101,8'b00000010,8'b00000100,8'b00000011,8'b11111111,8'b11011010,8'b00000100,8'b00000110,8'b11010110,8'b00000101,8'b11111100,8'b11111100,8'b00000111,8'b00000100,8'b00000001,8'b11010011,8'b00000011,8'b11111110,8'b11011001,8'b00000110,8'b00000011,8'b11110111,8'b00000100,8'b00000100,8'b00000001,8'b11011001,8'b11111100,8'b11111000,8'b11110011,8'b00001000,8'b00000100,8'b11101111,8'b00000010,8'b11111111,8'b00000001,8'b11100101,8'b11000111,8'b11100001,8'b00011100,8'b00011011,8'b00001000,8'b11110101,8'b00001101,8'b11011011,8'b00000001,8'b11111111,8'b00001001,8'b00001110,8'b11110100,8'b11011101,8'b11110101,8'b00011100,8'b11110111,8'b11001101,8'b11110110,8'b00000100,8'b00000110,8'b00010010,8'b11110001,8'b11110000,8'b11100001,8'b00010100,8'b11111010,8'b11001111,8'b11110011,8'b00000000,8'b00001000,8'b00001100,8'b11100100,8'b11111011,8'b11010010,8'b00001110,8'b11111001,8'b11110010,8'b11111010,8'b00000000,8'b00001000,8'b00001010,8'b11010100,8'b11111111,8'b11010100,8'b00001001,8'b00000001,8'b00000001,8'b11111110,8'b11101110,8'b00000101,8'b00000111,8'b11011010,8'b00000100,8'b11011100,8'b00000101,8'b00000010,8'b00000101,8'b00000001,8'b11001011,8'b11111111,8'b11111111,8'b11010000,8'b00000110,8'b11110100,8'b00000001,8'b00000001,8'b00000001,8'b00000101,8'b11010011,8'b11111110,8'b11111100,8'b11010101,8'b00001010,8'b00000001,8'b00000010,8'b00000100,8'b00000011,8'b00000111,8'b11100101,8'b11111001,8'b11101010,8'b11100110,8'b00010001,8'b00000111,8'b11110101,8'b00001000,8'b00000001,8'b00000101,8'b11101001,8'b11100010,8'b11000001,8'b00001110,8'b00011010,8'b00001000,8'b11100001,8'b00001010,8'b11101110,8'b11110011,8'b11101010,8'b00001110,8'b00010000,8'b11111001,8'b11100011,8'b11010101,8'b00100011,8'b11111110,8'b11011100,8'b11100000,8'b00000010,8'b00001000,8'b00001010,8'b11111000,8'b11111101,8'b11000101,8'b00010001,8'b00000101,8'b11100111,8'b11110010,8'b00000110,8'b00000110,8'b00000100,8'b11110111,8'b11111111,8'b10111111,8'b00001011,8'b00000111,8'b11111100,8'b11110101,8'b11111111,8'b00000001,8'b00000010,8'b11101100,8'b00000000,8'b11001100,8'b00001000,8'b00000001,8'b00000100,8'b11111011,8'b11101011,8'b11111100,8'b00000001,8'b11101100,8'b00000011,8'b11101100,8'b00000101,8'b11111110,8'b00000001,8'b00001011,8'b11010111,8'b11111111,8'b00000111,8'b11100011,8'b00001010,8'b11111110,8'b00001000,8'b00000010,8'b00000000,8'b00000111,8'b11010011,8'b11110010,8'b11111111,8'b11001110,8'b00001101,8'b00000100,8'b00000100,8'b11111110,8'b11110111,8'b00000100,8'b11110100,8'b11101101,8'b11110011,8'b11101011,8'b00001100,8'b00000010,8'b11110100,8'b00001000,8'b11110011,8'b11111100,8'b11111111,8'b11101111,8'b11100110,8'b00001010,8'b00010011,8'b11111011,8'b11101100,8'b00010110,8'b11011001,8'b11110010,8'b11111001,8'b11110000,8'b11111100,8'b00001111,8'b11110011,8'b11100110,8'b00010101,8'b11110101,8'b11110111,8'b11100000,8'b11111011,8'b11110111,8'b11111110,8'b00001101,8'b00000111,8'b11010110,8'b00000001,8'b00000110,8'b11111101,8'b11001111,8'b11111010,8'b11111100,8'b00000001,8'b00000111,8'b00000011,8'b11010001,8'b11111110,8'b00000010,8'b00001001,8'b11100101,8'b11110101,8'b11111111,8'b00000110,8'b00000111,8'b00000101,8'b11100001,8'b11111100,8'b00000100,8'b00001011,8'b11101110,8'b11101110,8'b11111011,8'b00000111,8'b00001011,8'b00000110,8'b00000010,8'b11110101,8'b11111101,8'b00001001,8'b11110110,8'b11001010,8'b11111001,8'b00001000,8'b00000000,8'b00001001,8'b00001001,8'b11111101,8'b00000001,8'b00000001,8'b11110111,8'b11001011,8'b11110010,8'b00001010,8'b11111111,8'b00001010,8'b00001101,8'b00000011,8'b00000111,8'b11101111,8'b11111100,8'b11101101,8'b11111011,8'b00000100,8'b11111111,8'b00000100,8'b00000101,8'b11111100,8'b00001000,8'b11011001,8'b11100001,8'b11111001,8'b00010101,8'b11101111,8'b00001111,8'b00000011,8'b00000011,8'b11111110,8'b00001111,8'b11010101,8'b11111011,8'b11111000,8'b11110100,8'b11111101,8'b00100000,8'b00000100,8'b11101111,8'b00001100,8'b11011111,8'b11111101,8'b11110100,8'b11111011,8'b11110111,8'b11111111,8'b00001101,8'b00001001,8'b11101101,8'b11111101,8'b11111100,8'b00000101,8'b11110000,8'b11110010,8'b11111010,8'b11111101,8'b00000111,8'b00000011,8'b11110011,8'b11111010,8'b11111010,8'b00000110,8'b11101101,8'b11101001,8'b00000010,8'b00000010,8'b00000111,8'b00000011,8'b11110100,8'b11111001,8'b11111110,8'b00001000,8'b11100110,8'b11010110,8'b11111111,8'b00000000,8'b00000011,8'b11111111,8'b11111011,8'b11101111,8'b11111010,8'b00000101,8'b11100110,8'b11011111,8'b00000000,8'b00001000,8'b00000001,8'b00000101,8'b00000100,8'b11111000,8'b00000100,8'b11111111,8'b11100100,8'b11011101,8'b00000010,8'b00000111,8'b00000111,8'b00000110,8'b00000111,8'b00001010,8'b00001001,8'b11101100,8'b11101100,8'b11110100,8'b00001011,8'b11111100,8'b00001100,8'b11111101,8'b00000011,8'b00001100,8'b00000100,8'b11011110,8'b11100000,8'b00001010,8'b00100101,8'b11011101,8'b00010011,8'b11011101,8'b11110011,8'b00000011,8'b11111000,8'b11100111,8'b11111110,8'b11111110,8'b00000110,8'b00001010,8'b00000111,8'b00000111,8'b11100101,8'b11111000,8'b11100000,8'b11101010,8'b00000001,8'b00001011,8'b11111101,8'b00000010,8'b00000001,8'b00000010,8'b11111110,8'b11111000,8'b11101110,8'b11111110,8'b11111110,8'b11111111,8'b11111101,8'b11111101,8'b11111111,8'b00000011,8'b11111100,8'b11111000,8'b11101111,8'b00000110,8'b11111111,8'b11110010,8'b11111101,8'b00000000,8'b00000100,8'b00000001,8'b00000000,8'b11111101,8'b11110100,8'b00000111,8'b00000100,8'b11110011,8'b00001001,8'b00001010,8'b00001010,8'b00000000,8'b00000110,8'b11111011,8'b11111110,8'b00000111,8'b00000000,8'b11111101,8'b00001010,8'b00000011,8'b11111111,8'b11111000,8'b00000100,8'b11111000,8'b11111100,8'b11110001,8'b00000100,8'b00000010,8'b00001111,8'b11111101,8'b00000101,8'b11110111,8'b00001010,8'b00001011,8'b11111111,8'b11011100,8'b00000111,8'b00001010,8'b00010001,8'b11101101,8'b00001011,8'b11100110,8'b00000100,8'b00001001,8'b11110100,8'b11011010,8'b00000010,8'b00010011,8'b00100000,8'b11001001,8'b00001001,8'b11000111,8'b11111111,8'b00000000,8'b11000100,8'b11100101,8'b00001001,8'b00011001,8'b00001000,8'b00001011,8'b11110110,8'b00000110,8'b11101111,8'b11101011,8'b11110101,8'b11100110,8'b00000001,8'b00001111,8'b00000001,8'b00001000,8'b11111000,8'b00000110,8'b11111100,8'b11101100,8'b00000000,8'b11110111,8'b11111111,8'b00000111,8'b00000001,8'b00000100,8'b11110111,8'b00000111,8'b00000000,8'b11101101,8'b00000001,8'b00000000,8'b00000011,8'b11111110,8'b00000011,8'b00000101,8'b11110101,8'b00000110,8'b00000110,8'b11101100,8'b00000110,8'b00000011,8'b00001000,8'b00000001,8'b00000110,8'b00001000,8'b11111000,8'b00000111,8'b00001001,8'b11101111,8'b00000110,8'b00000010,8'b00000011,8'b00000011,8'b00000011,8'b00000000,8'b11110001,8'b11111110,8'b00000111,8'b11101110,8'b00000000,8'b11110111,8'b11111110,8'b00000000,8'b00001000,8'b11111001,8'b11110101,8'b11110100,8'b00000000,8'b11101111,8'b11110111,8'b11101010,8'b11111110,8'b00001111,8'b00010010,8'b11110000,8'b00000100,8'b11101010,8'b00000010,8'b11110111,8'b11110100,8'b11111011,8'b11110010,8'b00001000,8'b00011110,8'b11011100,8'b11110111,8'b11010111,8'b11111100,8'b11101011,8'b11010110,8'b00001010,8'b00000010,8'b00010001,8'b00000011,8'b00001110,8'b11101001,8'b11111011,8'b10110100,8'b00001001,8'b11110000,8'b00001011,8'b00000000,8'b00000001,8'b11111101,8'b00001010,8'b11110011,8'b00000101,8'b11101100,8'b11111110,8'b00000001,8'b00000110,8'b11111111,8'b11111101,8'b11111111,8'b00000111,8'b11110000,8'b00000110,8'b11111010,8'b11111100,8'b00000011,8'b11111111,8'b11111111,8'b11111000,8'b11111011,8'b00000010,8'b11110001,8'b00000100,8'b11111011,8'b11110100,8'b00000000,8'b11111100,8'b00000110,8'b11111110,8'b00000010,8'b00001000,8'b11101111,8'b00000111,8'b00000101,8'b11110011,8'b00000111,8'b11111110,8'b00000011,8'b11111011,8'b11111111,8'b00000100,8'b11110010,8'b00000011,8'b00000100,8'b11101101,8'b00000001,8'b11111011,8'b11111101,8'b11111001,8'b11111101,8'b11110101,8'b11110100,8'b11111010,8'b11111010,8'b11100100,8'b11111110,8'b11111000,8'b11111000,8'b00000010,8'b00001011,8'b11111010,8'b00000011,8'b11111001,8'b11111010,8'b11011111,8'b00000000,8'b00000011,8'b11110011,8'b11111111,8'b00001000,8'b11011101,8'b00000110,8'b00000100,8'b11011001,8'b11011011,8'b11111111,8'b00010001,8'b11110101,8'b11111010,8'b00000011,8'b11111000,8'b11111101,8'b11110101,8'b00000101,8'b11110000,8'b11100010,8'b11011000,8'b11110011,8'b11111110,8'b00001100,8'b00001000,8'b11110001,8'b11110100,8'b00000111,8'b00000101,8'b11110011,8'b11000001,8'b11110001,8'b00001001,8'b00001011,8'b00000011,8'b11110000,8'b11110110,8'b11111100,8'b11110101,8'b11110000,8'b11100010,8'b11111010,8'b00001100,8'b00000010,8'b00001001,8'b00000011,8'b11111101,8'b00000010,8'b00000100,8'b11111100,8'b11010011,8'b11111100,8'b00000101,8'b11111010,8'b00000001,8'b11111010,8'b00001110,8'b00001001,8'b11011111,8'b11111010,8'b10101000,8'b00000110,8'b00001011,8'b11100011,8'b11110000,8'b00001011,8'b00001110,8'b00010110,8'b11000101,8'b11101101,8'b10000000,8'b11111110,8'b00101101,8'b10101010,8'b11010001,8'b00100101,8'b11100110,8'b00001010,8'b11101010,8'b00000000,8'b10101100,8'b11100111,8'b11111110,8'b11101100,8'b11110010,8'b00100111,8'b11111011,8'b00000011,8'b11000000,8'b00001101,8'b11000011,8'b11100000,8'b11110001,8'b11100101,8'b11111000,8'b11011100,8'b11111001,8'b00011111,8'b11011011,8'b00000000,8'b11110011,8'b11111110,8'b00000101,8'b00000011,8'b00000101,8'b00000011,8'b11111100,8'b11111111,8'b11111110,8'b11111011,8'b11111001,8'b11110000,8'b11101100,8'b11111111,8'b00000010,8'b11111011,8'b11111101,8'b11111011,8'b00000110,8'b11111101,8'b11110100,8'b11110011,8'b11111110,8'b00001001,8'b00000110,8'b00000010,8'b00000000,8'b11110110,8'b00010010,8'b11111101,8'b11111000,8'b11111001,8'b00000111,8'b00001001,8'b00000110,8'b11111110,8'b00000110,8'b00000000,8'b00001000,8'b00000011,8'b11110010,8'b00000011,8'b00001101,8'b11111110,8'b11111001,8'b00000010,8'b00000110,8'b00001011,8'b11011010,8'b11111001,8'b11011101,8'b11111010,8'b00100100,8'b11110000,8'b11101011,8'b00011101,8'b00000111,8'b00010000,8'b11100000,8'b11110100,8'b10111001,8'b11100001,8'b00011001,8'b10111010,8'b10111111,8'b00011110,8'b00001100,8'b00010001,8'b11011010,8'b00000010,8'b10111110,8'b11010100,8'b11110010,8'b10111100,8'b11011000,8'b00010111,8'b00011111,8'b00011101,8'b10110110,8'b00001011,8'b10101110,8'b11100000,8'b11111100,8'b11001010,8'b11011000,8'b00001000,8'b00001001,8'b00011100,8'b11010000,8'b11111100,8'b10110001,8'b11111110,8'b11110111,8'b00000011,8'b00000010,8'b11111111,8'b11111001,8'b11111010,8'b00000000,8'b00000001,8'b11111101,8'b11111000,8'b11101111,8'b11111111,8'b00000000,8'b11111011,8'b00000000,8'b11111010,8'b00000001,8'b00000000,8'b11111100,8'b11111100,8'b11100111,8'b00000011,8'b11111111,8'b11111110,8'b11111110,8'b11111011,8'b00000001,8'b00000010,8'b11111111,8'b00000000,8'b11111101,8'b00000011,8'b00000000,8'b11111010,8'b00000101,8'b00000001,8'b11110001,8'b00000011,8'b00001000,8'b11111101,8'b00010010,8'b11111110,8'b11111010,8'b00000011,8'b00000011,8'b00000110,8'b11100010,8'b11111000,8'b11110101,8'b11101110,8'b00010010,8'b00000101,8'b11100011,8'b00010100,8'b11111010,8'b00000100,8'b11100000,8'b11111011,8'b11110001,8'b11110011,8'b11111101,8'b11110110,8'b11101111,8'b00010100,8'b00010010,8'b00010000,8'b11100110,8'b11111011,8'b11110001,8'b11011110,8'b00000101,8'b11010001,8'b11110111,8'b00001011,8'b00011000,8'b00010001,8'b11110000,8'b11111111,8'b11011011,8'b11100110,8'b00001100,8'b11101001,8'b11110110,8'b00010111,8'b00001110,8'b00010001,8'b11110111,8'b11111101,8'b11010110,8'b00000010,8'b11111011,8'b11111010,8'b11110000,8'b11111011,8'b11110011,8'b11111111,8'b11111110,8'b11111010,8'b11111101,8'b00000101,8'b11101001,8'b11110110,8'b11111010,8'b00000110,8'b00000010,8'b00000011,8'b00000000,8'b00000111,8'b00000101,8'b11111110,8'b11101110,8'b11101111,8'b00000101,8'b00000010,8'b00000010,8'b11111111,8'b11111000,8'b11111011,8'b00000011,8'b11110010,8'b00000101,8'b11111000,8'b00010100,8'b11110000,8'b00000100,8'b11111100,8'b11100111,8'b11111010,8'b00000011,8'b11100111,8'b00010001,8'b00001010,8'b00001011,8'b11110110,8'b11100100,8'b11111000,8'b00001000,8'b11101011,8'b11111101,8'b00000110,8'b11100001,8'b00001000,8'b11101000,8'b00001110,8'b11101111,8'b00001010,8'b00000111,8'b11110101,8'b00000100,8'b00001110,8'b11111101,8'b00001001,8'b11111010,8'b11111101,8'b11111011,8'b11111111,8'b11111010,8'b00000000,8'b11110110,8'b11100111,8'b11111111,8'b11110100,8'b00000011,8'b00000100,8'b00000001,8'b11111100,8'b00000001,8'b00001001,8'b11110111,8'b11011011,8'b11111111,8'b11110111,8'b11111101,8'b00001001,8'b00000000,8'b11111110,8'b00000010,8'b00000111,8'b11110000,8'b00001011,8'b11111000,8'b00000101,8'b11110011,8'b00001011,8'b11111000,8'b00000101,8'b00000111,8'b11110111,8'b00000101,8'b00000100,8'b11101110,8'b11110101,8'b11111001,8'b00000101,8'b11111011,8'b00000001,8'b11110111,8'b11110001,8'b11111101,8'b11111100,8'b11111001,8'b11111000,8'b00010000,8'b11111111,8'b00000101,8'b00001000,8'b11110101,8'b11101111,8'b00000001,8'b11101011,8'b00000101,8'b11111110,8'b00100011,8'b11100111,8'b00000011,8'b00000000,8'b00000100,8'b11100110,8'b11101100,8'b11110101,8'b00010001,8'b11110111,8'b00010001,8'b11111011,8'b11101111,8'b11111101,8'b00010110,8'b11001011,8'b11111111,8'b00010000,8'b11110110,8'b00000000,8'b11110000,8'b00001101,8'b00000101,8'b00000000,8'b00011010,8'b11010011,8'b11111001,8'b00001011,8'b11111111,8'b00010000,8'b00000110,8'b11100011,8'b11101110,8'b11101100,8'b00000000,8'b00001100,8'b11111001,8'b11110110,8'b00000000,8'b00001101,8'b00001110,8'b00000101,8'b11001101,8'b11011011,8'b00000010,8'b00010011,8'b00000011,8'b11110100,8'b11111011,8'b00000111,8'b00000001,8'b00001111,8'b11011010,8'b11011110,8'b00000011,8'b00011010,8'b11111010,8'b00000010,8'b11100110,8'b00000010,8'b11110111,8'b00000011,8'b11111111,8'b11111100,8'b11111010,8'b11111001,8'b11110110,8'b00000010,8'b11101011,8'b00000111,8'b11101111,8'b11111111,8'b11110001,8'b11111110,8'b00000001,8'b11111100,8'b11110011,8'b00000011,8'b00000111,8'b00010010,8'b00000100,8'b11111010,8'b11110110,8'b00001111,8'b00010001,8'b00001000,8'b11110100,8'b11111001,8'b00010001,8'b00000100,8'b00001101,8'b11100111,8'b11111001,8'b00001111,8'b00001011,8'b11111011,8'b11011011,8'b00001000,8'b00010100,8'b11101001,8'b00000010,8'b11110101,8'b00000100,8'b00001101,8'b00010010,8'b11011111,8'b00000000,8'b00000011,8'b00001111,8'b11111110,8'b11111101,8'b11111100,8'b11111110,8'b11110011,8'b00001000,8'b11011110,8'b00000011,8'b11110101,8'b00000100,8'b00000101,8'b11111000,8'b00000101,8'b11010110,8'b11101011,8'b00000111,8'b00000100,8'b00001101,8'b00001001,8'b11101011,8'b00000110,8'b11111000,8'b00010010,8'b10111001,8'b11111110,8'b00001011,8'b00001010,8'b00000101,8'b00001011,8'b11110101,8'b00000101,8'b11011100,8'b00010011,8'b10111110,8'b00000111,8'b00000100,8'b00000101,8'b00000111,8'b00000001,8'b00000111,8'b00000111,8'b11111110,8'b00000001,8'b00000000,8'b11110001,8'b11110101,8'b00000101,8'b11101110,8'b11110110,8'b00000100,8'b00000000,8'b11111010,8'b11110010,8'b11111100,8'b11110101,8'b11110110,8'b00000011,8'b11101011,8'b11111101,8'b00000100,8'b00001010,8'b11111010,8'b11111000,8'b11111001,8'b00000010,8'b11111111,8'b00001000,8'b11110100,8'b11110011,8'b00001001,8'b00001011,8'b11110011,8'b11111000,8'b11101111,8'b00000011,8'b00000011,8'b00000100,8'b11111001,8'b11101100,8'b00010001,8'b11110100,8'b11110100,8'b00000000,8'b11101110,8'b11101110,8'b00000010,8'b11111001,8'b00000111,8'b11011110,8'b00011110,8'b00000011,8'b11101100,8'b00001101,8'b11110111,8'b11100100,8'b00001111,8'b11110000,8'b00010010,8'b00001100,8'b11101011,8'b11101111,8'b11111011,8'b00001010,8'b11110110,8'b00001011,8'b00001010,8'b11110011,8'b00001111,8'b00000100,8'b11000011,8'b11110101,8'b11111100,8'b00001101,8'b11101100,8'b00001100,8'b00011000,8'b11101011,8'b11111101,8'b00000101,8'b11110111,8'b11111111,8'b11101110,8'b00000010,8'b11100110,8'b00000111,8'b00010001,8'b11100001,8'b11111000,8'b11110110,8'b00001001,8'b00000010,8'b11111111,8'b11100111,8'b11110101,8'b11000111,8'b00001001,8'b11111100,8'b11110100,8'b11111010,8'b00001100,8'b00000100,8'b00000111,8'b00000001,8'b00001001,8'b11100011,8'b00000101,8'b00000110,8'b00000100,8'b11110100,8'b00000010,8'b00000011,8'b00000001,8'b00000010,8'b00001010,8'b11101010,8'b00000001,8'b11111110,8'b00000011,8'b11100100,8'b00001101,8'b00000001,8'b11111101,8'b00000100,8'b11111000,8'b11101000,8'b00000110,8'b11110111,8'b00000100,8'b11010110,8'b00010000,8'b00000001,8'b11101010,8'b00000111,8'b11111001,8'b11010011,8'b00001110,8'b11101100,8'b00001100,8'b00000001,8'b11110101,8'b11111000,8'b11111001,8'b00000011,8'b11111100,8'b11111100,8'b00001011,8'b11110111,8'b00001100,8'b00000101,8'b11011100,8'b11110010,8'b00001100,8'b11110011,8'b00000010,8'b00001000,8'b11111000,8'b11111110,8'b11111010,8'b11111110,8'b11101111,8'b11111101,8'b00001010,8'b11110011,8'b00000000,8'b00000101,8'b11111100,8'b11111110,8'b11110001,8'b00001110,8'b11111100,8'b00010010,8'b00001100,8'b11111100,8'b00000110,8'b00000111,8'b11110101,8'b00000000,8'b11110111,8'b11101110,8'b11110111,8'b11010101,8'b00011101,8'b00000110,8'b11110010,8'b11010000,8'b00001110,8'b11011100,8'b00001110,8'b11011001,8'b00000000,8'b11101000,8'b00010101,8'b00000111,8'b00000110,8'b10101000,8'b00010000,8'b11101011,8'b00001110,8'b10111000,8'b11111001,8'b11111100,8'b00001100,8'b00000100,8'b00001001,8'b10111101,8'b00001110,8'b11100011,8'b00001101,8'b11010100,8'b00000000,8'b11111101,8'b00000000,8'b00000100,8'b00000010,8'b11101111,8'b00001101,8'b11100000,8'b00001000,8'b11110011,8'b11111010,8'b11110111,8'b11111110,8'b00000000,8'b00000100,8'b11111010,8'b00000110,8'b11110100,8'b00000101,8'b00000010,8'b11111001,8'b11110101,8'b00001101,8'b11110111,8'b00000101,8'b11111111,8'b11111100,8'b00000100,8'b11111100,8'b00000000,8'b11111100,8'b11111100,8'b00000111,8'b11111001,8'b00000011,8'b00000010,8'b11110101,8'b00000100,8'b11110100,8'b11111011,8'b00000111,8'b00010000,8'b00000101,8'b11111010,8'b00000010,8'b11111011,8'b11101010,8'b00000011,8'b11101100,8'b00000000,8'b00000010,8'b00000001,8'b11111000,8'b00000010,8'b00000101,8'b11111000,8'b11101100,8'b00000010,8'b11111100,8'b11100000,8'b00001010,8'b11111010,8'b00000100,8'b11111000,8'b11101001,8'b00010100,8'b11101100,8'b11110011,8'b11111100,8'b11010110,8'b11111011,8'b00000001,8'b00000100,8'b11110001,8'b11011111,8'b00011111,8'b11101010,8'b11011000,8'b11011010,8'b11100100,8'b00001110,8'b00011110,8'b11111100,8'b11111000,8'b11100101,8'b00001100,8'b11100100,8'b11110011,8'b11001111,8'b11110000,8'b00001011,8'b00001111,8'b11111111,8'b00001011,8'b11101011,8'b00001111,8'b11100111,8'b11100010,8'b11000011,8'b11110110,8'b00001001,8'b00011010,8'b00001110,8'b11110001,8'b11100110,8'b00000110,8'b11010000,8'b00000100,8'b11110100,8'b11110100,8'b00001110,8'b00001100,8'b00000100,8'b11110110,8'b11101101,8'b00001000,8'b11001111,8'b11111101,8'b11101100,8'b11111001,8'b00001001,8'b00001110,8'b00000000,8'b11110100,8'b11111111,8'b00000101,8'b11011010,8'b00000111,8'b11010001,8'b11111101,8'b00001000,8'b00001010,8'b11111001,8'b11111100,8'b11111110,8'b00010001,8'b10110010,8'b00000100,8'b11011110,8'b11111001,8'b00000100,8'b00000010,8'b11100000,8'b00000110,8'b00000000,8'b00011001,8'b10111110,8'b11110100,8'b10110001,8'b11101100,8'b00010101,8'b11110000,8'b00000000,8'b00000111,8'b00000000,8'b00000000,8'b00000100,8'b11101111,8'b11010101,8'b11111100,8'b00000110,8'b11101100,8'b11101010,8'b00000111,8'b00000011,8'b00001001,8'b00000110,8'b00000011,8'b10111100,8'b00000100,8'b00011001,8'b11111100,8'b11111000,8'b00001101,8'b00001100,8'b00000110,8'b00000111,8'b11111110,8'b11010101,8'b11111010,8'b00010011,8'b11111100,8'b00000000,8'b00001001,8'b00000011,8'b11110110,8'b00000100,8'b11110011,8'b11011101,8'b00000001,8'b00001010,8'b00000110,8'b00001000,8'b00001100,8'b11111111,8'b11110111,8'b11111111,8'b11110100,8'b11101111,8'b00000110,8'b00001010,8'b00000111,8'b00000010,8'b00000101,8'b11101101,8'b11100010,8'b11111000,8'b11111100,8'b00000000,8'b00000111,8'b00000010,8'b00001010,8'b00000100,8'b00000101,8'b11100110,8'b11100000,8'b00000101,8'b00000100,8'b00001110,8'b00001100,8'b11111111,8'b00001000,8'b00000111,8'b11111110,8'b11110111,8'b11101011,8'b00000011,8'b00000111,8'b00000101,8'b00001100,8'b00001011,8'b00000011,8'b11111001,8'b00000000,8'b11111001,8'b11110011,8'b11111011,8'b00000001,8'b11110011,8'b11111011,8'b11110000,8'b11110011,8'b11111110,8'b00000110,8'b00000010,8'b00000010,8'b00000101,8'b11110000,8'b11101100,8'b11111110,8'b00000010,8'b11100100,8'b11110010,8'b00001010,8'b00000100,8'b00000101,8'b00000110,8'b11111110,8'b11110100,8'b11111011,8'b00000010,8'b11110111,8'b11110000,8'b00010010,8'b00001001,8'b00000010,8'b00010010,8'b00000100,8'b11101111,8'b11111001,8'b00010011,8'b11111000,8'b11111010,8'b00001110,8'b00000100,8'b11111000,8'b00001000,8'b00000110,8'b11100001,8'b11111101,8'b00000100,8'b00000011,8'b11111101,8'b00001001,8'b11110111,8'b11101001,8'b11111101,8'b11111100,8'b11111110,8'b00001000,8'b00000111,8'b00001100,8'b00000100,8'b00001011,8'b11100011,8'b11001010,8'b11111110,8'b00000110,8'b00000101,8'b00001111,8'b11101001,8'b00010001,8'b00001000,8'b00000110,8'b11001101,8'b11010100,8'b00000100,8'b00001010,8'b00001011,8'b00010001,8'b11100010,8'b00001011,8'b00000001,8'b11111010,8'b11011011,8'b11100101,8'b00001011,8'b00001111,8'b00001000,8'b00001011,8'b11111100,8'b11111101,8'b11110100,8'b11111011,8'b11100100,8'b11101111,8'b00000110,8'b00001010,8'b11111110,8'b00000011,8'b11111001,8'b11100111,8'b11100110,8'b00000101,8'b11111001,8'b00001111,8'b00001000,8'b00000001,8'b00000111,8'b00000001,8'b11111001,8'b11011011,8'b11011011,8'b00001000,8'b00000011,8'b00000100,8'b00000101,8'b00000101,8'b00000011,8'b11111100,8'b11110001,8'b11100110,8'b11100001,8'b00001111,8'b00001000,8'b00000101,8'b11111101,8'b00000111,8'b00000111,8'b11111001,8'b00001001,8'b11110001,8'b11110100,8'b00001100,8'b00000110,8'b11111111,8'b11101100,8'b00001101,8'b00001101,8'b11101000,8'b00000010,8'b11111000,8'b11110101,8'b11111100,8'b11110100,8'b11100111,8'b11110100,8'b00001000,8'b00000110,8'b00001101,8'b00000100,8'b00001011,8'b11110110,8'b00001011,8'b11110111,8'b11010011,8'b00000110,8'b00000010,8'b00000110,8'b00001011,8'b11100000,8'b00001001,8'b11110001,8'b00000000,8'b11110000,8'b11101000,8'b11111110,8'b11110111,8'b00000010,8'b00001110,8'b11110011,8'b00001010,8'b11110000,8'b00000001,8'b11110101,8'b11111011,8'b00000001,8'b11111100,8'b00000111,8'b00011000,8'b00010001,8'b00000111,8'b11010111,8'b11111001,8'b11011110,8'b00001110,8'b00000010,8'b11111011,8'b00001100,8'b00001001,8'b11111010,8'b11011100,8'b11100110,8'b00001001,8'b11101001,8'b00001011,8'b00001001,8'b00001001,8'b00001001,8'b00000110,8'b11111110,8'b11011010,8'b11100000,8'b00001001,8'b00000000,8'b00001000,8'b11111001,8'b00000110,8'b00001010,8'b00000001,8'b11011101,8'b11011110,8'b11110001,8'b00000111,8'b00000110,8'b00001011,8'b11101101,8'b00001001,8'b00000110,8'b11111100,8'b00000111,8'b11101001,8'b11110110,8'b00000011,8'b00000111,8'b00000011,8'b11101010,8'b00001101,8'b00001000,8'b11101100,8'b00000100,8'b11111001,8'b11111000,8'b11111010,8'b00000001,8'b11110110,8'b00000001,8'b00001011,8'b11111000,8'b00000011,8'b00000001,8'b00000000,8'b11110001,8'b00000110,8'b11111011,8'b11110001,8'b00001100,8'b11101001,8'b11111111,8'b00001010,8'b11110001,8'b11111111,8'b11111110,8'b00000000,8'b11111111,8'b11111100,8'b00000001,8'b11101000,8'b11110110,8'b00001110,8'b11101111,8'b11110100,8'b11111111,8'b11111100,8'b00000000,8'b00000010,8'b00000100,8'b11110101,8'b11111110,8'b00010000,8'b11011011,8'b11101100,8'b11111110,8'b11111110,8'b11111001,8'b00001000,8'b00000010,8'b11110100,8'b11111011,8'b00000100,8'b11010101,8'b00000001,8'b00000111,8'b00000101,8'b11110011,8'b11111110,8'b11111111,8'b11111001,8'b00001001,8'b00000111,8'b11010010,8'b11111101,8'b11111100,8'b00000100,8'b11111011,8'b00001011,8'b11110001,8'b00000100,8'b00000111,8'b00000111,8'b11110100,8'b11110101,8'b11111010,8'b11111100,8'b00000010,8'b00001001,8'b11100111,8'b00000011,8'b00000011,8'b11111011,8'b00000110,8'b11110101,8'b11111011,8'b11111001,8'b00000001,8'b00000101,8'b11101110,8'b00000110,8'b11111000,8'b11110111,8'b00000100,8'b11111010,8'b00000001,8'b11110101,8'b00000110,8'b11111101,8'b11111001,8'b11111111,8'b11101011,8'b11111110,8'b11111111,8'b11110101,8'b00000011,8'b00000001,8'b00000101,8'b00000000,8'b00000101,8'b11111010,8'b00000011,8'b00000111,8'b11110100,8'b11110000,8'b00000111,8'b11101111,8'b00000101,8'b00000101,8'b11111000,8'b00000011,8'b11111010,8'b00001010,8'b11111010,8'b11110000,8'b00000101,8'b11110010,8'b00000101,8'b00000101,8'b11111000,8'b00000100,8'b00000000,8'b00000001,8'b11101110,8'b11110101,8'b00000100,8'b11110110,8'b00000011,8'b11111101,8'b11110011,8'b00000110,8'b11111011,8'b00001000,8'b11011111,8'b00001000,8'b00001110,8'b11101110,8'b11111010,8'b11111001,8'b11101110,8'b11110111,8'b11110100,8'b00000111,8'b11100110,8'b00000100,8'b00000100,8'b11110001,8'b00000001,8'b00001000,8'b11100110,8'b00000000,8'b11111011,8'b00001001,8'b00000010,8'b00000101,8'b11111111,8'b11111000,8'b00000010,8'b00001010,8'b11101000,8'b00000100,8'b00000000,8'b00000110,8'b00000101,8'b11111110,8'b11111100,8'b11111000,8'b11111111,8'b00001000,8'b11110101,8'b00000010,8'b11110000,8'b11111101,8'b00001100,8'b11111010,8'b00000001,8'b11111100,8'b00000011,8'b00000110,8'b11111011,8'b00000010,8'b11111010,8'b11110101,8'b00000011,8'b11111010,8'b00000011,8'b00000101,8'b00000001,8'b00000000,8'b11111011,8'b00000100,8'b00000101,8'b11110000,8'b11110111,8'b11111000,8'b00000001,8'b11111011,8'b00000011,8'b11111101,8'b11101010,8'b00000110,8'b11111101,8'b11110011,8'b00001001,8'b11111011,8'b11111100,8'b11110010,8'b00000010,8'b11111101,8'b11100001,8'b00000011,8'b11111010,8'b11110100,8'b00000100,8'b11111001,8'b00000011,8'b11111111,8'b00001101,8'b11111001,8'b11101001,8'b00000000,8'b00001111,8'b00000100,8'b11110100,8'b00000110,8'b00010011,8'b11001111,8'b11111011,8'b11100000,8'b11101010,8'b00000100,8'b00000001,8'b00000101,8'b11111010,8'b00000100,8'b00001010,8'b11010111,8'b00000011,8'b11111100,8'b11011010,8'b00000110,8'b11111010,8'b00000100,8'b11111010,8'b00000010,8'b00000000,8'b11011110,8'b00000010,8'b00000001,8'b11101101,8'b00000010,8'b11111010,8'b00001110,8'b11111110,8'b00000000,8'b11111001,8'b11110010,8'b11111111,8'b00001100,8'b11111011,8'b00001011,8'b11111000,8'b00000100,8'b00001000,8'b11111001,8'b11110101,8'b00000001,8'b11111010,8'b00000101,8'b00000000,8'b00001001,8'b00000001,8'b11010111,8'b00000011,8'b00000100,8'b11111011,8'b00000111,8'b11111111,8'b11011011,8'b00000001,8'b00000101,8'b00000110,8'b11001110,8'b00000001,8'b00001000,8'b11111100,8'b00000101,8'b11110111,8'b11011100,8'b00000001,8'b00000011,8'b00000111,8'b11000100,8'b00010001,8'b00000101,8'b11110111,8'b00000100,8'b11111011,8'b11011111,8'b11110100,8'b11111100,8'b00000100,8'b11001011,8'b11111100,8'b11111101,8'b11100110,8'b00001000,8'b00000011,8'b11011010,8'b11101111,8'b11111111,8'b00010100,8'b11111100,8'b00001111,8'b11111110,8'b00011110,8'b11100011,8'b11110001,8'b11011100,8'b11110111,8'b00000011,8'b11101011,8'b11111110,8'b11111101,8'b11101110,8'b00010001,8'b11100101,8'b00000010,8'b10111101,8'b11111110,8'b00001000,8'b11111110,8'b00000100,8'b11111001,8'b11110011,8'b00001100,8'b11111011,8'b00001100,8'b11001010,8'b11111010,8'b00001010,8'b11111011,8'b00001110,8'b11111110,8'b11110110,8'b11111111,8'b11111100,8'b00000101,8'b11101111,8'b11111111,8'b00001001,8'b11111000,8'b11110110,8'b00000000,8'b11110101,8'b11011100,8'b00000100,8'b11110000,8'b11101100,8'b00001001,8'b00000010,8'b00000100,8'b10101010,8'b00010010,8'b11111110,8'b11100101,8'b00010000,8'b11100100,8'b11000100,8'b00001111,8'b11110011,8'b00001110,8'b10110100,8'b00011111,8'b00001011,8'b11101100,8'b00010011,8'b11011110,8'b11001001,8'b00001110,8'b11011011,8'b00001111,8'b11001100,8'b11111111,8'b00010100,8'b11010110,8'b11111111,8'b11110011,8'b11001011,8'b00001001,8'b11010010,8'b00010100,8'b11010011,8'b11100001,8'b11110000,8'b11110010,8'b00010001,8'b00000101,8'b11100100,8'b11111001,8'b11011010,8'b00010010,8'b11010101,8'b00111001,8'b00011011,8'b00001000,8'b11100011,8'b00010111,8'b11111111,8'b00001101,8'b11000110,8'b00000111};

	always_ff @(posedge clk) begin
		weight <= memory_B[weight_idx];  
   	end

	always_ff @(posedge clk) begin
		if ((mode != 1) && write_enable) 
            memory_A1[result_idx] <= result;

		data_a1 <= memory_A1[data_idx];
		
   	end
   	
	always_ff @(posedge clk) begin
		if ((mode == 1) && write_enable)
		        memory_A0[result_idx] <= result;

		data_a0 <= memory_A0[data_idx];
		
   	end
   	
   	//assign data_a1 = memory_A1[data_idx];
   	//assign data_a0 = memory_A0[data_idx];
   	assign data = (mode == 1) ? data_a1 : data_a0;

endmodule
